module domain

pub struct User {
	pub:
		user_id string
		display_name string
}