module redis

import domain { Event, Storage }

